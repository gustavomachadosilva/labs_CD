library verilog;
use verilog.vl_types.all;
entity E_dupla5 is
    port(
        S               : out    vl_logic;
        A               : in     vl_logic_vector(3 downto 0)
    );
end E_dupla5;
