library verilog;
use verilog.vl_types.all;
entity E_dupla5_vlg_vec_tst is
end E_dupla5_vlg_vec_tst;
