library verilog;
use verilog.vl_types.all;
entity ULA_BCD_vlg_vec_tst is
end ULA_BCD_vlg_vec_tst;
