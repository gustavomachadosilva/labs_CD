library verilog;
use verilog.vl_types.all;
entity COD_vlg_vec_tst is
end COD_vlg_vec_tst;
